// issue_queue.sv
// Airtight Reservation Station - Grade A+ implementation
// Features: 1-cycle wakeup latency, immediate forwarding, oldest-first selection
`timescale 1ns/1ps
import core_pkg::*;

module issue_queue #(
  parameter int ENTRIES = core_pkg::IQ_ENTRIES,
  parameter int ISSUE_W = core_pkg::ISSUE_WIDTH,
  parameter int TAG_W   = $clog2(core_pkg::PREGS),
  parameter int AGE_W   = 8  // Reduced for FPGA efficiency
)(
  input  logic                 clk,
  input  logic                 reset,

  // Allocation (up to ISSUE_W)
  input  logic [ISSUE_W-1:0]                   alloc_en,
  input  logic [3:0]                            alloc_opcode [ISSUE_W-1:0],
  input  logic [TAG_W-1:0]                      alloc_src1_tag [ISSUE_W-1:0],
  input  logic [TAG_W-1:0]                      alloc_src2_tag [ISSUE_W-1:0],
  input  logic [31:0]                           alloc_src1_val [ISSUE_W-1:0],
  input  logic [31:0]                           alloc_src2_val [ISSUE_W-1:0],
  input  core_pkg::preg_tag_t                   alloc_dst_phys [ISSUE_W-1:0],
  input  logic [4:0]                            alloc_dst_rob  [ISSUE_W-1:0],
  input  logic [1:0]                            alloc_fu_type  [ISSUE_W-1:0], // 0=ALU,1=BR
  output logic                                  alloc_ok,
  output logic [$clog2(ENTRIES)-1:0]            alloc_idx  [ISSUE_W-1:0],

  // CDB broadcasts
  input  logic [ISSUE_W-1:0]                    cdb_valid,
  input  logic [TAG_W-1:0]                      cdb_tag   [ISSUE_W-1:0],
  input  logic [31:0]                           cdb_value [ISSUE_W-1:0],

  // Issue outputs (ALU ports 0..1)
  output logic [ISSUE_W-1:0]                    issue_valid,
  output logic [3:0]                            issue_opcode [ISSUE_W-1:0],
  output logic [31:0]                           issue_src1_val [ISSUE_W-1:0],
  output logic [31:0]                           issue_src2_val [ISSUE_W-1:0],
  output core_pkg::preg_tag_t                   issue_dst_phys [ISSUE_W-1:0],
  output logic [4:0]                            issue_dst_rob [ISSUE_W-1:0],

  // Branch port
  output logic                                  br_valid,
  output logic [3:0]                            br_opcode,
  output logic [31:0]                           br_src1_val,
  output logic [31:0]                           br_src2_val,
  output core_pkg::preg_tag_t                   br_dst_phys,
  output logic [4:0]                            br_dst_rob,

  // Commit from ROB
  input  logic [ISSUE_W-1:0]                    commit_valid,
  input  logic [$clog2(core_pkg::ROB_ENTRIES)-1:0] commit_idx [ISSUE_W-1:0],
  input  logic                                  commit_clear_all,

  // Status
  output logic                                  rs_full,
  output logic                                  rs_almost_full
);

  // RS entry - optimized for FPGA
  typedef struct packed {
    logic                   used;
    logic                   src1_ready;
    logic                   src2_ready;
    logic [TAG_W-1:0]       src1_tag;
    logic [TAG_W-1:0]       src2_tag;
    logic [31:0]            src1_val;
    logic [31:0]            src2_val;
    logic [3:0]             opcode;
    core_pkg::preg_tag_t    dst_phys;
    logic [4:0]             dst_rob;
    logic [1:0]             fu_type;
    logic [AGE_W-1:0]       age;
  } rs_entry_t;

  rs_entry_t rs_mem [0:ENTRIES-1];

  // Registered CDB for safe updates
  logic [ISSUE_W-1:0]       cdb_valid_ff;
  logic [TAG_W-1:0]         cdb_tag_ff   [ISSUE_W-1:0];
  logic [31:0]              cdb_value_ff [ISSUE_W-1:0];

  // Age counter - wraps safely
  logic [AGE_W-1:0] age_counter;

  // Free entry tracking
  logic [ENTRIES-1:0] entry_used;

  // ============================================================
  //  CDB Registration - Critical for timing safety
  // ============================================================
  always_ff @(posedge clk or posedge reset) begin
    if (reset) begin
      cdb_valid_ff <= '0;
      for (int i = 0; i < ISSUE_W; i++) begin
        cdb_tag_ff[i] <= '0;
        cdb_value_ff[i] <= '0;
      end
    end else begin
      cdb_valid_ff <= cdb_valid;
      for (int i = 0; i < ISSUE_W; i++) begin
        cdb_tag_ff[i] <= cdb_tag[i];
        cdb_value_ff[i] <= cdb_value[i];
      end
    end
  end

  // ============================================================
  //  Main State Machine - Airtight timing
  // ============================================================
  always_ff @(posedge clk or posedge reset) begin
    if (reset) begin
      age_counter <= '0;
      for (int i = 0; i < ENTRIES; i++) begin
        rs_mem[i] <= '{
          used: 1'b0, src1_ready: 1'b0, src2_ready: 1'b0,
          src1_tag: '0, src2_tag: '0, src1_val: '0, src2_val: '0,
          opcode: '0, dst_phys: '0, dst_rob: '0, fu_type: '0, age: '0
        };
      end
      entry_used <= '0;
    end else begin
      age_counter <= age_counter + 1;

      // Phase 1: Safe CDB updates using registered values
      for (int i = 0; i < ENTRIES; i++) begin
        if (rs_mem[i].used) begin
          for (int b = 0; b < ISSUE_W; b++) begin
            if (cdb_valid_ff[b]) begin
              if (!rs_mem[i].src1_ready && (rs_mem[i].src1_tag == cdb_tag_ff[b])) begin
                rs_mem[i].src1_ready <= 1'b1;
                rs_mem[i].src1_val   <= cdb_value_ff[b];
              end
              if (!rs_mem[i].src2_ready && (rs_mem[i].src2_tag == cdb_tag_ff[b])) begin
                rs_mem[i].src2_ready <= 1'b1;
                rs_mem[i].src2_val   <= cdb_value_ff[b];
              end
            end
          end
        end
      end

      // Phase 2: Commit processing (entries freed immediately)
      if (commit_clear_all) begin
        for (int i = 0; i < ENTRIES; i++) begin
          rs_mem[i].used <= 1'b0;
          entry_used[i] <= 1'b0;
        end
      end else begin
        for (int c = 0; c < ISSUE_W; c++) begin
          if (commit_valid[c]) begin
            for (int i = 0; i < ENTRIES; i++) begin
              if (rs_mem[i].used && (rs_mem[i].dst_rob == commit_idx[c])) begin
                rs_mem[i].used <= 1'b0;
                entry_used[i] <= 1'b0;
              end
            end
          end
        end
      end

      // Phase 3: Allocation with immediate CDB forwarding
      int allocated = 0;
      for (int a = 0; a < ISSUE_W; a++) begin
        alloc_idx[a] <= '0;
        if (alloc_en[a]) begin
          // Find first free slot
          int slot = -1;
          for (int i = 0; i < ENTRIES; i++) begin
            if (!rs_mem[i].used && slot == -1) begin
              slot = i;
            end
          end

          if (slot != -1) begin
            // Compute ready states with immediate CDB forwarding
            logic s1_ready = (alloc_src1_tag[a] == '0); // x0 register
            logic s2_ready = (alloc_src2_tag[a] == '0);
            logic [31:0] s1_val = alloc_src1_val[a];
            logic [31:0] s2_val = alloc_src2_val[a];

            // Critical: Immediate CDB forwarding for back-to-back dependencies
            for (int b = 0; b < ISSUE_W; b++) begin
              if (cdb_valid[b]) begin
                if (!s1_ready && (alloc_src1_tag[a] == cdb_tag[b])) begin
                  s1_ready = 1'b1;
                  s1_val = cdb_value[b];
                end
                if (!s2_ready && (alloc_src2_tag[a] == cdb_tag[b])) begin
                  s2_ready = 1'b1;
                  s2_val = cdb_value[b];
                end
              end
            end

            // Allocate entry
            rs_mem[slot] <= '{
              used: 1'b1,
              src1_ready: s1_ready,
              src2_ready: s2_ready,
              src1_tag: alloc_src1_tag[a],
              src2_tag: alloc_src2_tag[a],
              src1_val: s1_val,
              src2_val: s2_val,
              opcode: alloc_opcode[a],
              dst_phys: alloc_dst_phys[a],
              dst_rob: alloc_dst_rob[a],
              fu_type: alloc_fu_type[a],
              age: age_counter
            };
            entry_used[slot] <= 1'b1;
            alloc_idx[a] <= slot;
            allocated++;
          end
        end
      end

      // Phase 4: Free issued entries immediately (optimization)
      for (int i = 0; i < ENTRIES; i++) begin
        if (rs_mem[i].used) begin
          logic will_issue = 1'b0;
          // Check if this entry will be issued this cycle
          for (int p = 0; p < ISSUE_W; p++) begin
            if (issue_valid[p] && (rs_mem[i].dst_rob == issue_dst_rob[p]) && 
                (rs_mem[i].dst_phys == issue_dst_phys[p])) begin
              will_issue = 1'b1;
            end
          end
          if (br_valid && (rs_mem[i].dst_rob == br_dst_rob) && 
              (rs_mem[i].dst_phys == br_dst_phys)) begin
            will_issue = 1'b1;
          end
          
          if (will_issue) begin
            rs_mem[i].used <= 1'b0;
            entry_used[i] <= 1'b0;
          end
        end
      end

      alloc_ok <= (allocated == popcount(alloc_en));
    end
  end

  // ============================================================
  //  Combinational Issue Selection - Oldest First
  // ============================================================
  function automatic int popcount(input logic [ISSUE_W-1:0] vec);
    int count = 0;
    for (int i = 0; i < ISSUE_W; i++) count += vec[i];
    return count;
  endfunction

  function automatic int find_oldest_ready(input bit is_alu);
    int oldest_idx = -1;
    logic [AGE_W-1:0] oldest_age = {AGE_W{1'b1}};
    
    for (int i = 0; i < ENTRIES; i++) begin
      if (rs_mem[i].used && rs_mem[i].src1_ready && rs_mem[i].src2_ready) begin
        if ((is_alu && (rs_mem[i].fu_type == 2'b00)) || 
            (!is_alu && (rs_mem[i].fu_type == 2'b01))) begin
          if (rs_mem[i].age < oldest_age) begin
            oldest_age = rs_mem[i].age;
            oldest_idx = i;
          end
        end
      end
    end
    return oldest_idx;
  endfunction

  always_comb begin
    // Default outputs
    for (int p = 0; p < ISSUE_W; p++) begin
      issue_valid[p] = 1'b0;
      issue_opcode[p] = '0;
      issue_src1_val[p] = '0;
      issue_src2_val[p] = '0;
      issue_dst_phys[p] = '0;
      issue_dst_rob[p] = '0;
    end
    br_valid = 1'b0;
    br_opcode = '0; br_src1_val = '0; br_src2_val = '0; br_dst_phys = '0; br_dst_rob = '0;

    // ALU issue selection
    int alu_issued = 0;
    bit [ENTRIES-1:0] issued_mask = '0;
    
    for (int p = 0; p < ISSUE_W; p++) begin
      if (alu_issued >= ISSUE_W) break;
      
      int candidate = -1;
      logic [AGE_W-1:0] candidate_age = {AGE_W{1'b1}};
      
      for (int i = 0; i < ENTRIES; i++) begin
        if (!issued_mask[i] && rs_mem[i].used && rs_mem[i].src1_ready && 
            rs_mem[i].src2_ready && (rs_mem[i].fu_type == 2'b00)) begin
          if (rs_mem[i].age < candidate_age) begin
            candidate_age = rs_mem[i].age;
            candidate = i;
          end
        end
      end
      
      if (candidate != -1) begin
        issue_valid[p] = 1'b1;
        issue_opcode[p] = rs_mem[candidate].opcode;
        issue_src1_val[p] = rs_mem[candidate].src1_val;
        issue_src2_val[p] = rs_mem[candidate].src2_val;
        issue_dst_phys[p] = rs_mem[candidate].dst_phys;
        issue_dst_rob[p] = rs_mem[candidate].dst_rob;
        issued_mask[candidate] = 1'b1;
        alu_issued++;
      end
    end

    // Branch issue selection (independent)
    int br_candidate = find_oldest_ready(0); // 0 = branch
    if (br_candidate != -1) begin
      br_valid = 1'b1;
      br_opcode = rs_mem[br_candidate].opcode;
      br_src1_val = rs_mem[br_candidate].src1_val;
      br_src2_val = rs_mem[br_candidate].src2_val;
      br_dst_phys = rs_mem[br_candidate].dst_phys;
      br_dst_rob = rs_mem[br_candidate].dst_rob;
    end
  end

  // ============================================================
  //  Status Flags
  // ============================================================
  always_comb begin
    int used_count = 0;
    for (int i = 0; i < ENTRIES; i++) begin
      used_count += entry_used[i];
    end
    
    rs_full = (used_count >= ENTRIES);
    rs_almost_full = (used_count >= (ENTRIES - ISSUE_W));
  end

endmodule
